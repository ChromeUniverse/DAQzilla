`default_nettype none

module top (
  // TODO: wire up modules
);

  // TODO: SPI core

  // TODO: DSP core

  // TODO: CAN core
  
endmodule